<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>13.3044,-73.3307,84.5552,-109.347</PageViewport>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-2,-12.5</position>
<gparam>LABEL_TEXT 1.Design 2X4 decoder using Cedar</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>12</ID>
<type>BA_DECODER_2x4</type>
<position>-10,-21</position>
<input>
<ID>ENABLE</ID>5 </input>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>5,-20</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>-16,-18.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>-19,-21.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>2.5,-16</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>8.5,-21.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>10.5,-24.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>-20.5,-24.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>BE_DECODER_3x8</type>
<position>-3,-32</position>
<input>
<ID>ENABLE</ID>8 </input>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>9 </input>
<output>
<ID>OUT_0</ID>19 </output>
<output>
<ID>OUT_1</ID>18 </output>
<output>
<ID>OUT_2</ID>17 </output>
<output>
<ID>OUT_3</ID>16 </output>
<output>
<ID>OUT_4</ID>15 </output>
<output>
<ID>OUT_5</ID>13 </output>
<output>
<ID>OUT_6</ID>12 </output>
<output>
<ID>OUT_7</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-14,-34.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>-8.5,-31.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-8,-37.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>-8,-28.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>18,-26</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>3.5,-29</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>11.5,-30</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>8,-31.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>5.5,-33</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>2,-34</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>12,-35</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>13.5,-37.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>BE_DECODER_3x8</type>
<position>2.5,-47.5</position>
<input>
<ID>ENABLE</ID>20 </input>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>22 </input>
<input>
<ID>IN_2</ID>21 </input>
<output>
<ID>OUT_1</ID>28 </output>
<output>
<ID>OUT_2</ID>29 </output>
<output>
<ID>OUT_3</ID>35 </output>
<output>
<ID>OUT_4</ID>30 </output>
<output>
<ID>OUT_5</ID>34 </output>
<output>
<ID>OUT_6</ID>33 </output>
<output>
<ID>OUT_7</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>-14,-40.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-45.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>-14.5,-49</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>-11.5,-53</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AE_OR4</type>
<position>27,-42.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>29 </input>
<input>
<ID>IN_3</ID>28 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_OR4</type>
<position>22,-52.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>35 </input>
<input>
<ID>IN_3</ID>32 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>53</ID>
<type>GA_LED</type>
<position>32,-42.5</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>27,-52.5</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>37.5,-42</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>32,-52</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,-16,1.5,-16</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-7,-19.5,-7,-16</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,-20,4,-20</points>
<connection>
<GID>14</GID>
<name>N_in0</name></connection>
<intersection>-7 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-7,-20.5,-7,-20</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,-21.5,7.5,-21.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<connection>
<GID>22</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-24.5,-7,-22.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-24.5,9.5,-24.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14,-18.5,-13,-18.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>-13 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13,-19.5,-13,-18.5</points>
<connection>
<GID>12</GID>
<name>ENABLE</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,-21.5,-13,-21.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,-24.5,-13,-22.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18.5,-24.5,-13,-24.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-28.5,-6,-28.5</points>
<connection>
<GID>28</GID>
<name>ENABLE</name></connection>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-33.5,-6,-31.5</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,-31.5,-6,-31.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-34.5,-6,-34.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-37.5,-6,-35.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-29,2.5,-29</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<intersection>0 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>0,-29.5,0,-29</points>
<connection>
<GID>28</GID>
<name>OUT_6</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-30,10.5,-30</points>
<connection>
<GID>37</GID>
<name>N_in0</name></connection>
<intersection>0 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>0,-30.5,0,-30</points>
<connection>
<GID>28</GID>
<name>OUT_5</name></connection>
<intersection>-30 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-28.5,0,-26</points>
<connection>
<GID>28</GID>
<name>OUT_7</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-26,17,-26</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>0,-31.5,7,-31.5</points>
<connection>
<GID>28</GID>
<name>OUT_4</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-33,4.5,-33</points>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<intersection>0 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>0,-33,0,-32.5</points>
<connection>
<GID>28</GID>
<name>OUT_3</name></connection>
<intersection>-33 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-34,0,-33.5</points>
<connection>
<GID>28</GID>
<name>OUT_2</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-34,1,-34</points>
<connection>
<GID>40</GID>
<name>N_in0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-35,11,-35</points>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<intersection>0 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>0,-35,0,-34.5</points>
<connection>
<GID>28</GID>
<name>OUT_1</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-37.5,0,-35.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-37.5,12.5,-37.5</points>
<connection>
<GID>42</GID>
<name>N_in0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-44,-0.5,-44</points>
<connection>
<GID>43</GID>
<name>ENABLE</name></connection>
<intersection>-12 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12,-44,-12,-40.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-49,-0.5,-49</points>
<connection>
<GID>43</GID>
<name>IN_2</name></connection>
<intersection>-11.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-11.5,-49,-11.5,-45.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-49 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-50,-5.5,-49</points>
<intersection>-50 2</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-49,-5.5,-49</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-50,-0.5,-50</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-53,-5.5,-51</points>
<intersection>-53 1</intersection>
<intersection>-51 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-53,-5.5,-53</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-51,-0.5,-51</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-50,14.5,-45.5</points>
<intersection>-50 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-45.5,24,-45.5</points>
<connection>
<GID>49</GID>
<name>IN_3</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-50,14.5,-50</points>
<connection>
<GID>43</GID>
<name>OUT_1</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-49,14.5,-43.5</points>
<intersection>-49 2</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-43.5,24,-43.5</points>
<connection>
<GID>49</GID>
<name>IN_2</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-49,14.5,-49</points>
<connection>
<GID>43</GID>
<name>OUT_2</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-47,14.5,-41.5</points>
<intersection>-47 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-41.5,24,-41.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-47,14.5,-47</points>
<connection>
<GID>43</GID>
<name>OUT_4</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-55.5,12.5,-39.5</points>
<intersection>-55.5 3</intersection>
<intersection>-44 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-39.5,24,-39.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-44,12.5,-44</points>
<connection>
<GID>43</GID>
<name>OUT_7</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>12.5,-55.5,19,-55.5</points>
<connection>
<GID>51</GID>
<name>IN_3</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-49.5,12,-45</points>
<intersection>-49.5 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-49.5,19,-49.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-45,12,-45</points>
<connection>
<GID>43</GID>
<name>OUT_6</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-51.5,12,-46</points>
<intersection>-51.5 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-51.5,19,-51.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-46,12,-46</points>
<connection>
<GID>43</GID>
<name>OUT_5</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-53.5,12,-48</points>
<intersection>-53.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-53.5,19,-53.5</points>
<connection>
<GID>51</GID>
<name>IN_2</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-48,12,-48</points>
<connection>
<GID>43</GID>
<name>OUT_3</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-42.5,31,-42.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<connection>
<GID>53</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-52.5,26,-52.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-18,39.1837,462.942,-203.926</PageViewport>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>48,-7.5</position>
<gparam>LABEL_TEXT 2.Design serial in and serial out shift resiter using D-ff</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AE_DFF_LOW_NT</type>
<position>-25,-17.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_DFF_LOW</type>
<position>10.5,-21</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clock</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_DFF_LOW</type>
<position>34.5,-21</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_DFF_LOW</type>
<position>71,-21.5</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>43 </output>
<input>
<ID>clock</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>-6,-19.5</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>75,-19.5</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>1,-15.5</position>
<gparam>LABEL_TEXT Data in</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>BB_CLOCK</type>
<position>-6.5,-24</position>
<output>
<ID>CLK</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>74,-15</position>
<gparam>LABEL_TEXT Data out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-19,31.5,-19</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>64</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-19.5,52.5,-19</points>
<intersection>-19.5 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-19.5,68,-19.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-19,52.5,-19</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,-19.5,7.5,-19.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>7.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7.5,-19.5,7.5,-19</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-19.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-26.5,68,-26.5</points>
<intersection>7.5 6</intersection>
<intersection>31.5 5</intersection>
<intersection>68 8</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>31.5,-26.5,31.5,-22</points>
<connection>
<GID>64</GID>
<name>clock</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>7.5,-26.5,7.5,-22</points>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<intersection>-26.5 1</intersection>
<intersection>-24 9</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>68,-26.5,68,-22.5</points>
<connection>
<GID>65</GID>
<name>clock</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-2.5,-24,7.5,-24</points>
<connection>
<GID>73</GID>
<name>CLK</name></connection>
<intersection>7.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-19.5,74,-19.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<connection>
<GID>70</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>118.769,-11.4854,270.942,-88.4069</PageViewport>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>59,12</position>
<gparam>LABEL_TEXT 2.Design serial in and serial out shift resiter using D-ff</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AE_DFF_LOW</type>
<position>21.5,-1.5</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>clock</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>77</ID>
<type>AE_DFF_LOW</type>
<position>45.5,-1.5</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>45 </output>
<input>
<ID>clock</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_DFF_LOW</type>
<position>82,-2</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_TOGGLE</type>
<position>5,0</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>86,0</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>12,4</position>
<gparam>LABEL_TEXT Data in</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>BB_CLOCK</type>
<position>4.5,-4.5</position>
<output>
<ID>CLK</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>85,4.5</position>
<gparam>LABEL_TEXT Data out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>32,7</position>
<input>
<ID>N_in2</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>GA_LED</type>
<position>62,7</position>
<input>
<ID>N_in2</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>60,-23.5</position>
<gparam>LABEL_TEXT 2.Design serial in and perallel out shift resiter using D-ff</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-37</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>54 </output>
<input>
<ID>clock</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_DFF_LOW</type>
<position>46.5,-37</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>55 </output>
<input>
<ID>clock</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_DFF_LOW</type>
<position>83,-37.5</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>clock</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_TOGGLE</type>
<position>6,-35.5</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>101</ID>
<type>GA_LED</type>
<position>87,-35.5</position>
<input>
<ID>N_in0</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>13,-31.5</position>
<gparam>LABEL_TEXT Data in</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>86,-31</position>
<gparam>LABEL_TEXT Data out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>GA_LED</type>
<position>33,-28.5</position>
<input>
<ID>N_in2</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>GA_LED</type>
<position>63,-28.5</position>
<input>
<ID>N_in2</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_TOGGLE</type>
<position>5,-41</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>173,12</position>
<gparam>LABEL_TEXT 3.Design perallell in and perallel out shift resiter using D-ff</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AE_DFF_LOW</type>
<position>135.5,-2</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>67 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>110</ID>
<type>AE_DFF_LOW</type>
<position>159.5,-2</position>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_DFF_LOW</type>
<position>196,-2.5</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>69 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_TOGGLE</type>
<position>131,4</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>113</ID>
<type>GA_LED</type>
<position>201.5,-11</position>
<input>
<ID>N_in3</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>119,-1.5</position>
<gparam>LABEL_TEXT Data in</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>199,4</position>
<gparam>LABEL_TEXT Data out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>140,-11.5</position>
<input>
<ID>N_in3</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>118,-6</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_TOGGLE</type>
<position>155,6</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_TOGGLE</type>
<position>190,5.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>121</ID>
<type>GA_LED</type>
<position>167,-11</position>
<input>
<ID>N_in3</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AE_DFF_LOW</type>
<position>144.5,-48</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>86 </output>
<input>
<ID>clock</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>123</ID>
<type>AE_DFF_LOW</type>
<position>164,-48</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>94 </output>
<input>
<ID>clock</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>124</ID>
<type>AE_DFF_LOW</type>
<position>204.5,-47</position>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>76 </output>
<input>
<ID>clock</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>126</ID>
<type>GA_LED</type>
<position>210,-55.5</position>
<input>
<ID>N_in3</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>132.5,-45</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>207.5,-40.5</position>
<gparam>LABEL_TEXT Serial out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>126,-51</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>172.5,-22.5</position>
<gparam>LABEL_TEXT 4.Design perallell in and seriel out shift resiter using D-ff</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_INVERTER</type>
<position>129.5,-28.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND2</type>
<position>146,-36.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_AND2</type>
<position>153.5,-36.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>164.5,-35.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>172,-35.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_TOGGLE</type>
<position>154.5,-25.5</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_OR2</type>
<position>149.5,-41.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_TOGGLE</type>
<position>173.5,-26</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>150</ID>
<type>AE_OR2</type>
<position>168.5,-40.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>136.5,-48</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>121,-28.5</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>150,-25.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AA_LABEL</type>
<position>170,-25.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>120.5,-24.5</position>
<gparam>LABEL_TEXT Load/shift</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,0.5,42.5,0.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>32 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>32,0.5,32,6</points>
<connection>
<GID>85</GID>
<name>N_in2</name></connection>
<intersection>0.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,0,63.5,0.5</points>
<intersection>0 1</intersection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,0,79,0</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,0.5,63.5,0.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>62 3</intersection>
<intersection>63.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>62,0.5,62,6</points>
<connection>
<GID>95</GID>
<name>N_in2</name></connection>
<intersection>0.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,0,18.5,0</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>18.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18.5,0,18.5,0.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>0 1</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-7,79,-7</points>
<intersection>18.5 6</intersection>
<intersection>42.5 5</intersection>
<intersection>79 8</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>42.5,-7,42.5,-2.5</points>
<connection>
<GID>77</GID>
<name>clock</name></connection>
<intersection>-7 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>18.5,-7,18.5,-2.5</points>
<connection>
<GID>76</GID>
<name>clock</name></connection>
<intersection>-7 1</intersection>
<intersection>-4.5 9</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>79,-7,79,-3</points>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>8.5,-4.5,18.5,-4.5</points>
<connection>
<GID>82</GID>
<name>CLK</name></connection>
<intersection>18.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,0,85,0</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<connection>
<GID>80</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-35,43.5,-35</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>33 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>33,-35,33,-29.5</points>
<connection>
<GID>105</GID>
<name>N_in2</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-35.5,64.5,-35</points>
<intersection>-35.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-35.5,80,-35.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-35,64.5,-35</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>63 3</intersection>
<intersection>64.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-35,63,-29.5</points>
<connection>
<GID>106</GID>
<name>N_in2</name></connection>
<intersection>-35 2</intersection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-35.5,19.5,-35.5</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19.5,-35.5,19.5,-35</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-42.5,80,-42.5</points>
<intersection>19.5 6</intersection>
<intersection>43.5 5</intersection>
<intersection>80 8</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43.5,-42.5,43.5,-38</points>
<connection>
<GID>98</GID>
<name>clock</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>19.5,-42.5,19.5,-38</points>
<connection>
<GID>97</GID>
<name>clock</name></connection>
<intersection>-42.5 1</intersection>
<intersection>-41 13</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>80,-42.5,80,-38.5</points>
<connection>
<GID>99</GID>
<name>clock</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>7,-41,19.5,-41</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>19.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-35.5,86,-35.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<connection>
<GID>101</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>132.5,-7.5,193,-7.5</points>
<intersection>132.5 6</intersection>
<intersection>156.5 5</intersection>
<intersection>193 8</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>156.5,-7.5,156.5,-3</points>
<connection>
<GID>110</GID>
<name>clock</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>132.5,-7.5,132.5,-3</points>
<connection>
<GID>109</GID>
<name>clock</name></connection>
<intersection>-7.5 1</intersection>
<intersection>-6 13</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>193,-7.5,193,-3.5</points>
<connection>
<GID>111</GID>
<name>clock</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>120,-6,132.5,-6</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>132.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,0,155,4</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155,0,156.5,0</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-0.5,190,3.5</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-0.5,193,-0.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,0,131,2</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,0,132.5,0</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-10.5,140,0</points>
<connection>
<GID>116</GID>
<name>N_in3</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,0,140,0</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-10,167,0</points>
<connection>
<GID>121</GID>
<name>N_in3</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,0,167,0</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-10,201.5,-0.5</points>
<connection>
<GID>113</GID>
<name>N_in3</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199,-0.5,201.5,-0.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>201.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128.5,-53,201.5,-53</points>
<intersection>128.5 30</intersection>
<intersection>141.5 31</intersection>
<intersection>159.5 5</intersection>
<intersection>201.5 8</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>159.5,-53,159.5,-49</points>
<intersection>-53 1</intersection>
<intersection>-49 34</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>201.5,-53,201.5,-48</points>
<connection>
<GID>124</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>128.5,-53,128.5,-51</points>
<intersection>-53 1</intersection>
<intersection>-51 39</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>141.5,-53,141.5,-49</points>
<connection>
<GID>122</GID>
<name>clock</name></connection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>34</ID>
<points>159.5,-49,161,-49</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>159.5 5</intersection></hsegment>
<hsegment>
<ID>39</ID>
<points>128,-51,128.5,-51</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>128.5 30</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-54.5,210,-45</points>
<connection>
<GID>126</GID>
<name>N_in3</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207.5,-45,210,-45</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>132.5,-28.5,171,-28.5</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>152.5 8</intersection>
<intersection>171 9</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>152.5,-33.5,152.5,-28.5</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>171,-32.5,171,-28.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-33.5,154.5,-27.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126.5,-31,165.5,-31</points>
<intersection>126.5 2</intersection>
<intersection>147 4</intersection>
<intersection>165.5 5</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126.5,-31,126.5,-28.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-31 1</intersection>
<intersection>-28.5 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>147,-33.5,147,-31</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-31 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>165.5,-32.5,165.5,-31</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>123,-28.5,126.5,-28.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>126.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-39,148.5,-38.5</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>-39 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>146,-39.5,146,-39</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>146,-39,148.5,-39</points>
<intersection>146 1</intersection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-39.5,153.5,-39</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<intersection>-39 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>150.5,-39,150.5,-38.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>150.5,-39,153.5,-39</points>
<intersection>150.5 1</intersection>
<intersection>153.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-42.5,141,-33.5</points>
<intersection>-42.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-42.5,147.5,-42.5</points>
<intersection>141 0</intersection>
<intersection>147.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-33.5,145,-33.5</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>141 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>147.5,-46,147.5,-42.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>149.5,-46,161,-46</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>149.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>149.5,-46,149.5,-44.5</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-32.5,173,-30</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-30 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>173.5,-30,173.5,-28</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>173,-30,173.5,-30</points>
<intersection>173 0</intersection>
<intersection>173.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>164.5,-38.5,164.5,-38</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>164.5,-38,167.5,-38</points>
<intersection>164.5 1</intersection>
<intersection>167.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>167.5,-38,167.5,-37.5</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-38 2</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>172,-38.5,172,-37.5</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>169.5,-37.5,172,-37.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>172 1</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-44,168.5,-43.5</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168.5,-44,201.5,-44</points>
<intersection>168.5 0</intersection>
<intersection>201.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>201.5,-45,201.5,-44</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-43,160,-32.5</points>
<intersection>-43 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-43,167,-43</points>
<intersection>160 0</intersection>
<intersection>167 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,-32.5,163.5,-32.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>167,-46,167,-43</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>-43 1</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>141.5,-48,141.5,-46</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-48 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>138.5,-48,141.5,-48</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>141.5 4</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-61.7877,7.87753,208.742,-128.872</PageViewport>
<gate>
<ID>4</ID>
<type>BB_CLOCK</type>
<position>14.5,-34.5</position>
<output>
<ID>CLK</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BE_JKFF_LOW</type>
<position>27.5,-26.5</position>
<input>
<ID>J</ID>25 </input>
<input>
<ID>K</ID>25 </input>
<output>
<ID>Q</ID>31 </output>
<input>
<ID>clock</ID>24 </input>
<output>
<ID>nQ</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7</ID>
<type>BE_JKFF_LOW</type>
<position>72.5,-25.5</position>
<input>
<ID>J</ID>26 </input>
<input>
<ID>K</ID>26 </input>
<output>
<ID>Q</ID>36 </output>
<input>
<ID>clock</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>11.5,-26.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>63.5,-18.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>15</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>100.5,-26.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>36 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>17</ID>
<type>BB_CLOCK</type>
<position>14,-66.5</position>
<output>
<ID>CLK</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 2</lparam></gate>
<gate>
<ID>19</ID>
<type>BE_JKFF_LOW</type>
<position>27,-58.5</position>
<input>
<ID>J</ID>50 </input>
<input>
<ID>K</ID>50 </input>
<output>
<ID>Q</ID>63 </output>
<input>
<ID>clock</ID>49 </input>
<output>
<ID>nQ</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>21</ID>
<type>BE_JKFF_LOW</type>
<position>72.5,-57.5</position>
<input>
<ID>J</ID>51 </input>
<input>
<ID>K</ID>51 </input>
<output>
<ID>Q</ID>71 </output>
<input>
<ID>clock</ID>52 </input>
<output>
<ID>nQ</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>11,-58.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>63,-50.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>100,-58.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>71 </input>
<input>
<ID>IN_2</ID>73 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>58,-46</position>
<gparam>LABEL_TEXT 5.Design 3 bit asycro counter using positive adge trigger and t-ff</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>BE_JKFF_LOW</type>
<position>91,-56</position>
<input>
<ID>J</ID>60 </input>
<input>
<ID>K</ID>60 </input>
<output>
<ID>Q</ID>73 </output>
<input>
<ID>clock</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>83,-49</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>BB_CLOCK</type>
<position>11,-99</position>
<output>
<ID>CLK</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 2</lparam></gate>
<gate>
<ID>55</ID>
<type>BE_JKFF_LOW</type>
<position>24,-91</position>
<input>
<ID>J</ID>75 </input>
<input>
<ID>K</ID>75 </input>
<output>
<ID>Q</ID>88 </output>
<input>
<ID>clock</ID>74 </input>
<output>
<ID>nQ</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>58</ID>
<type>BE_JKFF_LOW</type>
<position>69.5,-90</position>
<input>
<ID>J</ID>78 </input>
<input>
<ID>K</ID>78 </input>
<output>
<ID>Q</ID>93 </output>
<input>
<ID>clock</ID>79 </input>
<output>
<ID>nQ</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>8,-91</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>60,-83</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>66</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>152,-104</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>93 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>98 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>55,-78.5</position>
<gparam>LABEL_TEXT 6.Design 3 bit asycro counter using positive adge trigger and t-ff</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>BE_JKFF_LOW</type>
<position>88.5,-88.5</position>
<input>
<ID>J</ID>80 </input>
<input>
<ID>K</ID>80 </input>
<output>
<ID>Q</ID>96 </output>
<input>
<ID>clock</ID>81 </input>
<output>
<ID>nQ</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>80.5,-81.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>84</ID>
<type>BE_JKFF_LOW</type>
<position>131,-84.5</position>
<input>
<ID>J</ID>100 </input>
<input>
<ID>K</ID>100 </input>
<output>
<ID>Q</ID>98 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>124,-68.5</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>58.5,-14</position>
<gparam>LABEL_TEXT 4.Design 2 bit asycro counter using positive adge trigger and t-ff</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-34.5,21.5,-26.5</points>
<intersection>-34.5 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-26.5,24.5,-26.5</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-34.5,21.5,-34.5</points>
<connection>
<GID>4</GID>
<name>CLK</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-28.5,17,-24.5</points>
<intersection>-28.5 1</intersection>
<intersection>-26.5 3</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-28.5,24.5,-28.5</points>
<connection>
<GID>6</GID>
<name>K</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-24.5,24.5,-24.5</points>
<connection>
<GID>6</GID>
<name>J</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>13.5,-26.5,17,-26.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-27.5,63.5,-20.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-27.5,69.5,-27.5</points>
<connection>
<GID>7</GID>
<name>K</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-23.5,69.5,-23.5</points>
<connection>
<GID>7</GID>
<name>J</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-28.5,50,-25.5</points>
<intersection>-28.5 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-25.5,69.5,-25.5</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-28.5,50,-28.5</points>
<connection>
<GID>6</GID>
<name>nQ</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-31.5,97.5,-31.5</points>
<intersection>30.5 3</intersection>
<intersection>97.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,-31.5,30.5,-24.5</points>
<connection>
<GID>6</GID>
<name>Q</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>97.5,-31.5,97.5,-27.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-26.5,86.5,-23.5</points>
<intersection>-26.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-26.5,97.5,-26.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-23.5,86.5,-23.5</points>
<connection>
<GID>7</GID>
<name>Q</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-66.5,21,-58.5</points>
<intersection>-66.5 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-58.5,24,-58.5</points>
<connection>
<GID>19</GID>
<name>clock</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-66.5,21,-66.5</points>
<connection>
<GID>17</GID>
<name>CLK</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-60.5,16.5,-56.5</points>
<intersection>-60.5 1</intersection>
<intersection>-58.5 3</intersection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-60.5,24,-60.5</points>
<connection>
<GID>19</GID>
<name>K</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-56.5,24,-56.5</points>
<connection>
<GID>19</GID>
<name>J</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>13,-58.5,16.5,-58.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-59.5,63,-52.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-59.5 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-59.5,69.5,-59.5</points>
<connection>
<GID>21</GID>
<name>K</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-55.5,69.5,-55.5</points>
<connection>
<GID>21</GID>
<name>J</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-60.5,49.5,-57.5</points>
<intersection>-60.5 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-57.5,69.5,-57.5</points>
<connection>
<GID>21</GID>
<name>clock</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-60.5,49.5,-60.5</points>
<connection>
<GID>19</GID>
<name>nQ</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-58,83,-51</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-58 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-58,88,-58</points>
<connection>
<GID>34</GID>
<name>K</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,-54,88,-54</points>
<connection>
<GID>34</GID>
<name>J</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-59.5,81,-56</points>
<intersection>-59.5 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-56,88,-56</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-59.5,81,-59.5</points>
<connection>
<GID>21</GID>
<name>nQ</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-68.5,95,-68.5</points>
<intersection>30 3</intersection>
<intersection>95 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30,-68.5,30,-56.5</points>
<connection>
<GID>19</GID>
<name>Q</name></connection>
<intersection>-68.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>95,-68.5,95,-59.5</points>
<intersection>-68.5 1</intersection>
<intersection>-59.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>95,-59.5,97,-59.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>95 4</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-64,97,-64</points>
<intersection>75.5 3</intersection>
<intersection>97 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75.5,-64,75.5,-55.5</points>
<connection>
<GID>21</GID>
<name>Q</name></connection>
<intersection>-64 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>97,-64,97,-58.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-64 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-57.5,95.5,-54</points>
<intersection>-57.5 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-57.5,97,-57.5</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,-54,95.5,-54</points>
<connection>
<GID>34</GID>
<name>Q</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-99,18,-91</points>
<intersection>-99 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-91,21,-91</points>
<connection>
<GID>55</GID>
<name>clock</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-99,18,-99</points>
<connection>
<GID>52</GID>
<name>CLK</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-93,13.5,-89</points>
<intersection>-93 1</intersection>
<intersection>-91 3</intersection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-93,21,-93</points>
<connection>
<GID>55</GID>
<name>K</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-89,21,-89</points>
<connection>
<GID>55</GID>
<name>J</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>10,-91,13.5,-91</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-92,60,-85</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>-92 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-92,66.5,-92</points>
<connection>
<GID>58</GID>
<name>K</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-88,66.5,-88</points>
<connection>
<GID>58</GID>
<name>J</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-93,46.5,-90</points>
<intersection>-93 2</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-90,66.5,-90</points>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-93,46.5,-93</points>
<connection>
<GID>55</GID>
<name>nQ</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-90.5,80.5,-83.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-90.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-90.5,85.5,-90.5</points>
<connection>
<GID>69</GID>
<name>K</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-86.5,85.5,-86.5</points>
<connection>
<GID>69</GID>
<name>J</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-92,78,-88.5</points>
<intersection>-92 2</intersection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-88.5,85.5,-88.5</points>
<connection>
<GID>69</GID>
<name>clock</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-92,78,-92</points>
<connection>
<GID>58</GID>
<name>nQ</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-101,97,-101</points>
<intersection>27 3</intersection>
<intersection>97 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-101,27,-89</points>
<connection>
<GID>55</GID>
<name>Q</name></connection>
<intersection>-101 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>97,-105,97,-101</points>
<intersection>-105 5</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>97,-105,149,-105</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>97 4</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-96.5,94,-96.5</points>
<intersection>72.5 3</intersection>
<intersection>94 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72.5,-96.5,72.5,-88</points>
<connection>
<GID>58</GID>
<name>Q</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>94,-104,94,-96.5</points>
<intersection>-104 7</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>94,-104,149,-104</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>94 4</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-103,92.5,-86.5</points>
<intersection>-103 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-103,149,-103</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-86.5,92.5,-86.5</points>
<connection>
<GID>69</GID>
<name>Q</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-102,142,-82.5</points>
<intersection>-102 1</intersection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-102,149,-102</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134,-82.5,142,-82.5</points>
<connection>
<GID>84</GID>
<name>Q</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-90.5,109.5,-84.5</points>
<intersection>-90.5 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-84.5,128,-84.5</points>
<connection>
<GID>84</GID>
<name>clock</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-90.5,109.5,-90.5</points>
<connection>
<GID>69</GID>
<name>nQ</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-86.5,121,-82.5</points>
<intersection>-86.5 2</intersection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-82.5,128,-82.5</points>
<connection>
<GID>84</GID>
<name>J</name></connection>
<intersection>121 0</intersection>
<intersection>124 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-86.5,128,-86.5</points>
<connection>
<GID>84</GID>
<name>K</name></connection>
<intersection>121 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>124,-82.5,124,-70.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-82.5 1</intersection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>75.6872,22.2452,237.504,-59.5514</PageViewport>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>144.5,-8.5</position>
<gparam>LABEL_TEXT 6. 2 bit asychronous up down</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>BE_JKFF_LOW</type>
<position>120.5,-22.5</position>
<input>
<ID>J</ID>101 </input>
<input>
<ID>K</ID>101 </input>
<output>
<ID>Q</ID>114 </output>
<input>
<ID>clock</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>91</ID>
<type>BE_JKFF_LOW</type>
<position>149.5,-23.5</position>
<input>
<ID>J</ID>107 </input>
<input>
<ID>K</ID>107 </input>
<output>
<ID>Q</ID>113 </output>
<input>
<ID>clock</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>107.5,-23.5</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>129,-36.5</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>117</ID>
<type>AO_XNOR2</type>
<position>128.5,-30.5</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>171.5,-23</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>113 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>141</ID>
<type>BB_CLOCK</type>
<position>107.5,-34</position>
<output>
<ID>CLK</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_TOGGLE</type>
<position>140.5,-31</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>148.5,-38</position>
<gparam>LABEL_TEXT 0 up</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>149,-43.5</position>
<gparam>LABEL_TEXT 1 down</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>132.5,-40</position>
<gparam>LABEL_TEXT Modifire</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-24.5,113,-20.5</points>
<intersection>-24.5 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-24.5,117.5,-24.5</points>
<connection>
<GID>90</GID>
<name>K</name></connection>
<intersection>109.5 5</intersection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113,-20.5,117.5,-20.5</points>
<connection>
<GID>90</GID>
<name>J</name></connection>
<intersection>113 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>109.5,-24.5,109.5,-23.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129,-33.5,129.5,-33.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-34.5,129,-33.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-25.5,140,-21.5</points>
<intersection>-25.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,-25.5,146.5,-25.5</points>
<connection>
<GID>91</GID>
<name>K</name></connection>
<intersection>140 0</intersection>
<intersection>140.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,-21.5,146.5,-21.5</points>
<connection>
<GID>91</GID>
<name>J</name></connection>
<intersection>140 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>140.5,-29,140.5,-25.5</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-27.5,128.5,-23.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-23.5,146.5,-23.5</points>
<connection>
<GID>91</GID>
<name>clock</name></connection>
<intersection>128.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-34,114.5,-22.5</points>
<intersection>-34 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-22.5,117.5,-22.5</points>
<connection>
<GID>90</GID>
<name>clock</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-34,114.5,-34</points>
<connection>
<GID>141</GID>
<name>CLK</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,-23,160.5,-21.5</points>
<intersection>-23 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160.5,-23,168.5,-23</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>152.5,-21.5,160.5,-21.5</points>
<connection>
<GID>91</GID>
<name>Q</name></connection>
<intersection>160.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-19,146,-18.5</points>
<intersection>-19 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146,-19,165.5,-19</points>
<intersection>146 0</intersection>
<intersection>165.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-18.5,146,-18.5</points>
<intersection>125.5 3</intersection>
<intersection>146 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>125.5,-33.5,125.5,-18.5</points>
<intersection>-33.5 7</intersection>
<intersection>-20.5 6</intersection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>165.5,-24,165.5,-19</points>
<intersection>-24 5</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>165.5,-24,168.5,-24</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>165.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>123.5,-20.5,125.5,-20.5</points>
<connection>
<GID>90</GID>
<name>Q</name></connection>
<intersection>125.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>125.5,-33.5,127.5,-33.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>125.5 3</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>76.7128,12.5626,228.886,-64.3589</PageViewport>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>132.5,-3.5</position>
<gparam>LABEL_TEXT 7. Sycronous counter with sequence 0,1,3,5,7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>BE_JKFF_LOW</type>
<position>108,-25.5</position>
<input>
<ID>J</ID>116 </input>
<output>
<ID>Q</ID>117 </output>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>165</ID>
<type>BE_JKFF_LOW</type>
<position>124,-25</position>
<input>
<ID>clock</ID>115 </input>
<output>
<ID>nQ</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>166</ID>
<type>BE_JKFF_LOW</type>
<position>148.5,-24.5</position>
<input>
<ID>clock</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>168</ID>
<type>BB_CLOCK</type>
<position>95.5,-31.5</position>
<output>
<ID>CLK</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>170</ID>
<type>GA_LED</type>
<position>112.5,-11</position>
<input>
<ID>N_in2</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-34.5,102,-31.5</points>
<intersection>-34.5 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-34.5,141.5,-34.5</points>
<intersection>102 0</intersection>
<intersection>105 5</intersection>
<intersection>118 3</intersection>
<intersection>141.5 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99.5,-31.5,102,-31.5</points>
<connection>
<GID>168</GID>
<name>CLK</name></connection>
<intersection>102 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>118,-34.5,118,-25</points>
<intersection>-34.5 1</intersection>
<intersection>-25 8</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>105,-34.5,105,-25.5</points>
<connection>
<GID>164</GID>
<name>clock</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>141.5,-34.5,141.5,-24.5</points>
<intersection>-34.5 1</intersection>
<intersection>-24.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>141.5,-24.5,145.5,-24.5</points>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<intersection>141.5 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>118,-25,121,-25</points>
<connection>
<GID>165</GID>
<name>clock</name></connection>
<intersection>118 3</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-17.5,129,-17.5</points>
<intersection>105 4</intersection>
<intersection>129 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>129,-27,129,-17.5</points>
<intersection>-27 5</intersection>
<intersection>-17.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>105,-23.5,105,-17.5</points>
<connection>
<GID>164</GID>
<name>J</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>127,-27,129,-27</points>
<connection>
<GID>165</GID>
<name>nQ</name></connection>
<intersection>129 3</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-23.5,112.5,-12</points>
<connection>
<GID>170</GID>
<name>N_in2</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-23.5,112.5,-23.5</points>
<connection>
<GID>164</GID>
<name>Q</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>0,39.1837,480.942,-203.926</PageViewport></page 6>
<page 7>
<PageViewport>0,39.1837,480.942,-203.926</PageViewport></page 7>
<page 8>
<PageViewport>0,39.1837,480.942,-203.926</PageViewport></page 8>
<page 9>
<PageViewport>0,39.1837,480.942,-203.926</PageViewport></page 9></circuit>